/home/mingliu/bluedbm/src/lib/AuroraGearbox.bsv